module basic_layer_search(

);

Ref_mem Ref_mem();

PE_array PE_array();

SAD_Tree SAD_Tree();

endmodule